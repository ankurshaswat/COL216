library IEEE;
use IEEE.std_logic_1164.all;


entity Main_Controller is
  port (
    ins_20 : in std_logic;
    ins_31_28 : in std_logic_vector(3 downto 0);
    ins_27_26 : in std_logic_vector(1 downto 0);
    F         : in std_logic_vector(3 downto 0);  -- (Flags : Z & N & V & C )
    p         : in std_logic;
    clk       : in std_logic;
--CONTROL SIGNALS
    --------------

    IorD  : out std_logic;
--MR: out std_logic:='0';
    MW    : out std_logic;
    IW    : out std_logic;
    DW    : out std_logic;
    Rsrc  : out std_logic;
    M2R   : out std_logic_vector(1 downto 0);  --
    RW    : out std_logic;
    AW    : out std_logic;
    BW    : out std_logic;
    Asrc1 : out std_logic_vector(1 downto 0);  --
    Asrc2 : out std_logic_vector(1 downto 0);
    Fset  : out std_logic;
    op    : out std_logic_vector(3 downto 0);
    ReW   : out std_logic;

    WadSrc      : out std_logic_vector(1 downto 0);
    R1src       : out std_logic_vector(1 downto 0);
    op1sel      : out std_logic;
    SType       : out std_logic_vector(1 downto 0);
    ShiftAmtSel : out std_logic;
    Shift       : out std_logic;
    MulW        : out std_logic;
    ShiftW      : out std_logic;
    op1update   : out std_logic
    );
end entity Main_Controller;

architecture arch of Main_Controller is

  type state_type is (fetch, rdAB, arith, addr, brn, wrRF, wrM, rdM, M2RF, shift_state, readx, rdM_and_auto_incr_res2RF, wrMRF, addr_rdB);
  signal state : state_type;

  signal Z, N, V, C : std_logic;

begin

  process (clk)
  begin
    if (rising_edge(clk)) then
      case state is

--------------------------------------------|        
		when fetch =>
          IorD  <= '0';
          --MR: out std_logic:='0';
          --  PW          <= '1';
          MW    <= '0';
          IW    <= '1';
          DW    <= '0';
          Rsrc  <= '0';
          M2R   <= "00";                --
          RW    <= '0';
          AW    <= '0';
          BW    <= '0';
          Asrc1 <= "00";
          Asrc2 <= "01";
          Fset  <= '0';
          op    <= "0100";
          ReW   <= '0';

          WadSrc      <= "000";
          R1src       <= "00";
          op1sel      <= '0';
          SType       <= "00";
          ShiftAmtSel <= '0';
          Shift       <= '0';
          MulW        <= '0';
          ShiftW      <= '0';
          op1update   <= '0';
          state       <= rdAB;
--------------------------------------------|
        when rdAB =>

          if (ins_27_26 = "00") then
            state <= arith;
            IorD  <= '0';
            --MR: out std_logic:='0';
            --  PW          <= '0';
            MW    <= '0';
            IW    <= '0';
            DW    <= '0';
            Rsrc  <= '0';
            M2R   <= "00";              --
            RW    <= '0';
            AW    <= '1';
            BW    <= '1';
            Asrc1 <= "00";
            Asrc2 <= "01";
            Fset  <= '0';
            op    <= "0100";
            ReW   <= '0';

            WadSrc      <= "000";
            R1src       <= "01";
            op1sel      <= '0';
            SType       <= "00";
            ShiftAmtSel <= '0';
            Shift       <= '0';
            MulW        <= '0';
            ShiftW      <= '0';
            op1update   <= '0';
          elsif (ins_27_26 = "01") then state <= addr;
          elsif (ins_27_26 = "10") then state <= brn;
          end if;
--------------------------------------------|
        when arith =>
          state <= wrRF;
--------------------------------------------|
        when addr =>
          if (ins_20 = '0') then state <= wrM;
          else state                   <= rdM;
          end if;
--------------------------------------------|
        when wrM =>
          state <= fetch;
--------------------------------------------|
        when rdM =>
          state <= M2RF;
--------------------------------------------|
        when brn =>
          state <= fetch;
--------------------------------------------|
        when wrRF =>
          state <= fetch;
--------------------------------------------|
        when M2RF =>
          state <= fetch;
--------------------------------------------|
        when shift_state =>
          if (ins_27_26 = "00") then state   <= arith;
          elsif(ins_27_26 = "01") then state <= addr_rdB;
          end if;
--------------------------------------------|
        when readx =>
          state <= shift_state;
--------------------------------------------|
        when rdM_and_auto_incr_res2RF =>
          if (ins_20 = '0') then state <= wrMRF;
          else state                   <= M2RF;
          end if;
--------------------------------------------|
        when  wrMRF =>
            state <= fetch;
--------------------------------------------|
        when  addr_rdB =>
            state <= rdM_and_auto_incr_res2RF;


      end case;
    end if;
  end process;



end architecture;
